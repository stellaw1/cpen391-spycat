
//////////////////////////////////////////////////////////////////////////////////
// Top level WHOLE system not just Qsys generated HPS system
//////////////////////////////////////////////////////////////////////////////////

module spycat (
		/////////////////////////////////////////////
		// FPGA Pins
		/////////////////////////////////////////////
	
		// Clock pins
		input CLOCK_50,CLOCK2_50,CLOCK3_50,CLOCK4_50, 
		
		// Seven Segment Displays
		// These are the names of the 6 seven segment display on the DE1 and those in the PIN Planner,
		//	so stick to these names.
		output unsigned [6:0] HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,
	
		// Pushbuttons
		input unsigned [3:0] KEY,
	
		// LEDs
		output unsigned [9:0] LEDR,
	
		// Slider Switches
		input unsigned [9:0] SW,
		
		// VGA/Graphics Signals
		output VGA_BLANK_N,
		output VGA_SYNC_N,
		output VGA_CLK,
		output VGA_HS,
		output VGA_VS,
		
		output unsigned [7:0] VGA_B,
		output unsigned [7:0] VGA_G,
		output unsigned [7:0] VGA_R,
	
		// SDRAM on FPGA Side
		output unsigned [12:0] DRAM_ADDR,
		output unsigned [1:0] DRAM_BA,
		output DRAM_CAS_N,
		output DRAM_CKE,
		output DRAM_CLK,
		output DRAM_CS_N,
		inout unsigned [15:0] DRAM_DQ,
		output DRAM_LDQM,
		output DRAM_RAS_N,
		output DRAM_UDQM,
		output DRAM_WE_N,
		
		// 40-Pin Headers
		inout unsigned [35:0] GPIO_0,
		inout unsigned [35:0] GPIO_1,
		

		//////////////////////////////////////////////////////
		// HPS Pins
		//////////////////////////////////////////////////////
		
		// DDR3 SDRAM
		output unsigned [14:0] HPS_DDR3_ADDR,
		output unsigned [2:0] HPS_DDR3_BA,
		output HPS_DDR3_CAS_N,
		output HPS_DDR3_CKE,
		output HPS_DDR3_CK_N,
		output HPS_DDR3_CK_P,
		output HPS_DDR3_CS_N,
		output unsigned [3:0] HPS_DDR3_DM,
		inout unsigned [31:0] HPS_DDR3_DQ,
		inout unsigned [3:0] HPS_DDR3_DQS_N,
		inout unsigned [3:0] HPS_DDR3_DQS_P,
		output HPS_DDR3_ODT,
		output HPS_DDR3_RAS_N,
		output HPS_DDR3_RESET_N	,
		input HPS_DDR3_RZQ,
		output HPS_DDR3_WE_N,
		
		// Ethernet
		output HPS_ENET_GTX_CLK,
		inout HPS_ENET_INT_N,
		output HPS_ENET_MDC,
		inout HPS_ENET_MDIO,
		input HPS_ENET_RX_CLK,
		input unsigned [3:0] HPS_ENET_RX_DATA,
		input HPS_ENET_RX_DV,
		output unsigned [3:0] HPS_ENET_TX_DATA,
		output HPS_ENET_TX_EN,
	
		// Flash
		inout unsigned [3:0] HPS_FLASH_DATA,
		output HPS_FLASH_DCLK,
		output HPS_FLASH_NCSO,
	
		// Accelerometer
		inout HPS_GSENSOR_INT,
			
		// General Purpose I/O
		inout unsigned [1:0] HPS_GPIO,
		
		// I2C
		inout HPS_I2C_CONTROL,
		inout HPS_I2C1_SCLK,
		inout HPS_I2C1_SDAT,
		inout HPS_I2C2_SCLK,
		inout HPS_I2C2_SDAT,
	
		// Pushbutton
		inout HPS_KEY,
	
		// LED
		inout HPS_LED,
			
		// SD Card
		output HPS_SD_CLK,
		inout HPS_SD_CMD,
		inout unsigned [3:0] HPS_SD_DATA,
	
		// SPI
		output HPS_SPIM_CLK,
		input HPS_SPIM_MISO,
		output HPS_SPIM_MOSI,
		inout HPS_SPIM_SS,
	
		// UART
		input HPS_UART_RX,
		output HPS_UART_TX,
	
		// USB
		inout HPS_CONV_USB_N,
		input HPS_USB_CLKOUT,
		inout unsigned [7:0] HPS_USB_DATA,
		input HPS_USB_DIR,
		input HPS_USB_NXT,
		output HPS_USB_STP 
	 );

///////////////////////////////////////////////////////////////////////////////////////////
//  signal declarations for temporary signals/wires to connect sub-systems together
///////////////////////////////////////////////////////////////////////////////////////////

	 // temp wires carrying 2 sets of 4 bit data to each pair of Hex displays
	 // The 3 pairs of 8 bit ports generated by QSYS will drive these wires
	 // and they will be connected to the 7-Segment decoders created in VHDL 
	 // and they will drive the real HEX display on the DE1
	 
	 wire unsigned [7:0] Temp_hex0_1;
	 wire unsigned [7:0] Temp_hex2_3;
	 wire unsigned [7:0] Temp_hex4_5;

	 wire unsigned [1:0] Temp_SDRAM_DQM;
	 
	 
	// TEMP Wires  TO CONNECT IO BRIDGE from QSYS generated IOBridge TO SUBSYSTEMS INCLUDING GRAPHICS AND IO DEVICE (RS232'S)
   
	reg IO_ACK_WIRE;									// reg because driven by always@ block
	wire IO_IRQ_WIRE;
	wire unsigned [15:0] IO_Address_WIRE;
	wire IO_Bus_Enable_WIRE;
	wire unsigned [1:0] IO_Byte_Enable_WIRE;
	wire IO_RW_WIRE;
	wire unsigned [15:0] IO_Write_Data_WIRE;
	wire unsigned [15:0] IO_Read_Data_WIRE;

	// camera
	// wire unsigned [9:0] MIPI_pixel_D;
	// wire MIPI_refclk;
	// wire MIPI_reset;
	// wire MIPI_pixel_clk;
	// wire MIPI_pixel_HS;
	// wire MIPI_pixel_VS;
	// wire MIPI_chip_select;
	// wire MIPI_I2C_scl;
	// wire MIPI_I2C_sda;
	// wire MIPI_mclk;
	// wire camera_pwdwn;
	// wire camera_I2C_scl;
	// wire camera_I2C_sda;

	wire unsigned [28:0] hps_sdram_address;
	wire unsigned [7:0] hps_sdram_burstcount;	
	wire hps_sdram_waitrequest;	
	wire unsigned [31:0] hps_sdram_writedata;	
	wire hps_sdram_write;

	wire unsigned [31:0] hps_sdram_readdata;
	wire hps_sdram_readdatavalid;
	wire hps_sdram_read;

	wire [31:0] cmd_from_hps;
	wire unsigned [28:0] camera_out_address;	
	wire unsigned [25:0] camera_out_data;	
	wire camera_out_write, camera_fps;
	
	// Other temporary wires 
	wire RESET_L_WIRE;
	wire IO_Enable_L_WIRE;
	wire IO_UpperByte_Select_L_WIRE;
	wire IO_LowerByte_Select_L_WIRE;
	
	// for LCD display connected to PIO port, 11 bits used
	wire unsigned [15:0] LCD_WIRE;
 
	 ///////////////////////////////////////////////////////////////////////////////////////
	 // u0 is an instanace of the QSYS generated computer
	 // map its IO ports as described below
	 ///////////////////////////////////////////////////////////////////////////////////////
	 
		 CPEN391_Computer u0 (
//			.hex0_1_export                   (Temp_hex0_1),                   //               hex0_1.export
//			.hex2_3_export                   (Temp_hex2_3),                   //               hex2_3.export
//			.hex4_5_export                   (Temp_hex4_5),                   //               hex4_5.export
			.hps_io_hps_io_emac1_inst_TX_CLK (HPS_ENET_GTX_CLK), 					//               hps_io.hps_io_emac1_inst_TX_CLK
			.hps_io_hps_io_emac1_inst_TXD0   (HPS_ENET_TX_DATA[0]),   			//                     .hps_io_emac1_inst_TXD0
			.hps_io_hps_io_emac1_inst_TXD1   (HPS_ENET_TX_DATA[1]),   			//                     .hps_io_emac1_inst_TXD1
			.hps_io_hps_io_emac1_inst_TXD2   (HPS_ENET_TX_DATA[2]),   			//                     .hps_io_emac1_inst_TXD2
			.hps_io_hps_io_emac1_inst_TXD3   (HPS_ENET_TX_DATA[3]),   			//                     .hps_io_emac1_inst_TXD3
			.hps_io_hps_io_emac1_inst_RXD0   (HPS_ENET_RX_DATA[0]),   			//                     .hps_io_emac1_inst_RXD0
			.hps_io_hps_io_emac1_inst_MDIO   (HPS_ENET_MDIO),   					//                     .hps_io_emac1_inst_MDIO
			.hps_io_hps_io_emac1_inst_MDC    (HPS_ENET_MDC),    					//                     .hps_io_emac1_inst_MDC
			.hps_io_hps_io_emac1_inst_RX_CTL (HPS_ENET_RX_DV), 					//                     .hps_io_emac1_inst_RX_CTL
			.hps_io_hps_io_emac1_inst_TX_CTL (HPS_ENET_TX_EN), 					//                     .hps_io_emac1_inst_TX_CTL
			.hps_io_hps_io_emac1_inst_RX_CLK (HPS_ENET_RX_CLK), 					//                     .hps_io_emac1_inst_RX_CLK
			.hps_io_hps_io_emac1_inst_RXD1   (HPS_ENET_RX_DATA[1]),   			//                     .hps_io_emac1_inst_RXD1
			.hps_io_hps_io_emac1_inst_RXD2   (HPS_ENET_RX_DATA[2]),   			//                     .hps_io_emac1_inst_RXD2
			.hps_io_hps_io_emac1_inst_RXD3   (HPS_ENET_RX_DATA[3]),   			//                     .hps_io_emac1_inst_RXD3
			.hps_io_hps_io_qspi_inst_IO0     (HPS_FLASH_DATA[0]),     			//                     .hps_io_qspi_inst_IO0
			.hps_io_hps_io_qspi_inst_IO1     (HPS_FLASH_DATA[1]),     			//                     .hps_io_qspi_inst_IO1
			.hps_io_hps_io_qspi_inst_IO2     (HPS_FLASH_DATA[2]),     			//                     .hps_io_qspi_inst_IO2
			.hps_io_hps_io_qspi_inst_IO3     (HPS_FLASH_DATA[3]),     			//                     .hps_io_qspi_inst_IO3
			.hps_io_hps_io_qspi_inst_SS0     (HPS_FLASH_NCSO),     				//                     .hps_io_qspi_inst_SS0
			.hps_io_hps_io_qspi_inst_CLK     (HPS_FLASH_DCLK),     				//                     .hps_io_qspi_inst_CLK
			.hps_io_hps_io_sdio_inst_CMD     (HPS_SD_CMD),     					//                     .hps_io_sdio_inst_CMD
			.hps_io_hps_io_sdio_inst_D0      (HPS_SD_DATA[0]),      				//                     .hps_io_sdio_inst_D0
			.hps_io_hps_io_sdio_inst_D1      (HPS_SD_DATA[1]),      				//                     .hps_io_sdio_inst_D1
			.hps_io_hps_io_sdio_inst_CLK     (HPS_SD_CLK),     					//                     .hps_io_sdio_inst_CLK
			.hps_io_hps_io_sdio_inst_D2      (HPS_SD_DATA[2]),      				//                     .hps_io_sdio_inst_D2
			.hps_io_hps_io_sdio_inst_D3      (HPS_SD_DATA[3]),      				//                     .hps_io_sdio_inst_D3
			.hps_io_hps_io_usb1_inst_D0      (HPS_USB_DATA[0]),      			//                     .hps_io_usb1_inst_D0
			.hps_io_hps_io_usb1_inst_D1      (HPS_USB_DATA[1]),      			//                     .hps_io_usb1_inst_D1
			.hps_io_hps_io_usb1_inst_D2      (HPS_USB_DATA[2]),      			//                     .hps_io_usb1_inst_D2
			.hps_io_hps_io_usb1_inst_D3      (HPS_USB_DATA[3]),      			//                     .hps_io_usb1_inst_D3
			.hps_io_hps_io_usb1_inst_D4      (HPS_USB_DATA[4]),      			//                     .hps_io_usb1_inst_D4
			.hps_io_hps_io_usb1_inst_D5      (HPS_USB_DATA[5]),      			//                     .hps_io_usb1_inst_D5
			.hps_io_hps_io_usb1_inst_D6      (HPS_USB_DATA[6]),      			//                     .hps_io_usb1_inst_D6
			.hps_io_hps_io_usb1_inst_D7      (HPS_USB_DATA[7]),      			//                     .hps_io_usb1_inst_D7
			.hps_io_hps_io_usb1_inst_CLK     (HPS_USB_CLKOUT),     				//                     .hps_io_usb1_inst_CLK
			.hps_io_hps_io_usb1_inst_STP     (HPS_USB_STP),     					//                     .hps_io_usb1_inst_STP
			.hps_io_hps_io_usb1_inst_DIR     (HPS_USB_DIR),     					//                     .hps_io_usb1_inst_DIR
			.hps_io_hps_io_usb1_inst_NXT     (HPS_USB_NXT),     					//                     .hps_io_usb1_inst_NXT
			.hps_io_hps_io_spim1_inst_CLK    (HPS_SPIM_CLK),    					//                     .hps_io_spim1_inst_CLK
			.hps_io_hps_io_spim1_inst_MOSI   (HPS_SPIM_MOSI),   					//                     .hps_io_spim1_inst_MOSI
			.hps_io_hps_io_spim1_inst_MISO   (HPS_SPIM_MISO),   					//                     .hps_io_spim1_inst_MISO
			.hps_io_hps_io_spim1_inst_SS0    (HPS_SPIM_SS),    					//                     .hps_io_spim1_inst_SS0
			.hps_io_hps_io_uart0_inst_RX     (HPS_UART_RX),     					//                     .hps_io_uart0_inst_RX
			.hps_io_hps_io_uart0_inst_TX     (HPS_UART_TX),     					//                     .hps_io_uart0_inst_TX
			.hps_io_hps_io_i2c0_inst_SDA     (HPS_I2C1_SDAT),     				//                     .hps_io_i2c0_inst_SDA
			.hps_io_hps_io_i2c0_inst_SCL     (HPS_I2C1_SCLK),     				//                     .hps_io_i2c0_inst_SCL
			.hps_io_hps_io_i2c1_inst_SDA     (HPS_I2C2_SDAT),     				//                     .hps_io_i2c1_inst_SDA
			.hps_io_hps_io_i2c1_inst_SCL     (HPS_I2C2_SCLK),     				//                     .hps_io_i2c1_inst_SCL
			.hps_io_hps_io_gpio_inst_GPIO09  (HPS_CONV_USB_N),  					//                     .hps_io_gpio_inst_GPIO09
			.hps_io_hps_io_gpio_inst_GPIO35  (HPS_ENET_INT_N),  					//                     .hps_io_gpio_inst_GPIO35
			.hps_io_hps_io_gpio_inst_GPIO40  (HPS_GPIO[0]),  						//                     .hps_io_gpio_inst_GPIO40
			.hps_io_hps_io_gpio_inst_GPIO41  (HPS_GPIO[1]),  						//                     .hps_io_gpio_inst_GPIO41
			.hps_io_hps_io_gpio_inst_GPIO48  (HPS_I2C_CONTROL),  					//                     .hps_io_gpio_inst_GPIO48
			.hps_io_hps_io_gpio_inst_GPIO53  (HPS_LED),  							//                     .hps_io_gpio_inst_GPIO53
			.hps_io_hps_io_gpio_inst_GPIO54  (HPS_KEY),  							//                     .hps_io_gpio_inst_GPIO54
			.hps_io_hps_io_gpio_inst_GPIO61  (HPS_GSENSOR_INT),  					//                     .hps_io_gpio_inst_GPIO61

			// IO Bridge Connections to wires
			.io_acknowledge  						(IO_ACK_WIRE),	
			.io_irq          						(IO_IRQ_WIRE),
			.io_address      						(IO_Address_WIRE),
			.io_bus_enable  						(IO_Bus_Enable_WIRE),
			.io_byte_enable  						(IO_Byte_Enable_WIRE),
			.io_rw           						(IO_RW_WIRE),  
			.io_write_data   						(IO_Write_Data_WIRE),                    
			.io_read_data    						(IO_Read_Data_WIRE),

			// 2x24 LCD Display Connections to 16 bit PIO port
			// .lcd_export								(LCD_WIRE),

			
			// Red LED connections
			//!!!.leds_export                     (LEDR),                     		//                 leds.export
			
			// SDRAM connections on the FPGA side
			.memory_mem_a                    (HPS_DDR3_ADDR),                 //               memory.mem_a
			.memory_mem_ba                   (HPS_DDR3_BA),                   //                     .mem_ba
			.memory_mem_ck                   (HPS_DDR3_CK_P),                 //                     .mem_ck
			.memory_mem_ck_n                 (HPS_DDR3_CK_N),                 //                     .mem_ck_n
			.memory_mem_cke                  (HPS_DDR3_CKE),                  //                     .mem_cke
			.memory_mem_cs_n                 (HPS_DDR3_CS_N),                 //                     .mem_cs_n
			.memory_mem_ras_n                (HPS_DDR3_RAS_N),                //                     .mem_ras_n
			.memory_mem_cas_n                (HPS_DDR3_CAS_N),                //                     .mem_cas_n
			.memory_mem_we_n                 (HPS_DDR3_WE_N),                 //                     .mem_we_n
			.memory_mem_reset_n              (HPS_DDR3_RESET_N),              //                     .mem_reset_n
			.memory_mem_dq                   (HPS_DDR3_DQ),                   //                     .mem_dq
			.memory_mem_dqs                  (HPS_DDR3_DQS_P),                //                     .mem_dqs
			.memory_mem_dqs_n                (HPS_DDR3_DQS_N),                //                     .mem_dqs_n
			.memory_mem_odt                  (HPS_DDR3_ODT),                  //                     .mem_odt
			.memory_mem_dm                   (HPS_DDR3_DM),                   //                     .mem_dm
			.memory_oct_rzqin                (HPS_DDR3_RZQ),                	//                     .oct_rzqin
//			.pushbuttons_export              (KEY),              					//          pushbuttons.export
			.sdram_pll_refclk_clk 			 (CLOCK_50),
			.new_sdram_controller_0_addr	 (DRAM_ADDR),  // new_sdram_controller_0_wire.addr
			.new_sdram_controller_0_ba	 	 (DRAM_BA),    //                            .ba
			.new_sdram_controller_0_cas_n	 (DRAM_CAS_N), //                            .cas_n
			.new_sdram_controller_0_cke	 	 (DRAM_CKE),   //                            .cke
			.new_sdram_controller_0_cs_n	 (DRAM_CS_N),  //                            .cs_n
			.new_sdram_controller_0_dq	 	 (DRAM_DQ),    //                            .dq
			.new_sdram_controller_0_dqm	 	 ({DRAM_UDQM, DRAM_LDQM}),   //                            .dqm
			.new_sdram_controller_0_ras_n	 (DRAM_RAS_N), //                            .ras_n
			.new_sdram_controller_0_we_n	 (DRAM_WE_N),  // 
			.sdram_clk_1_clk                 (DRAM_CLK),                   	//            sdram_clk.clk
			// .sdram_addr                      (DRAM_ADDR),                     //                sdram.addr
			// .sdram_ba                        (DRAM_BA),                       //                     .ba
			// .sdram_cas_n                     (DRAM_CAS_N),                    //                     .cas_n
			// .sdram_cke                       (DRAM_CKE),                      //                     .cke
			// .sdram_cs_n                      (DRAM_CS_N),                     //                     .cs_n
			// .sdram_dq                        (DRAM_DQ),                       //                     .dq
			// .sdram_dqm 		                (Temp_SDRAM_DQM),                //                     .dqm
			// .sdram_ras_n                     (DRAM_RAS_N),                    //                     .ras_n
			// .sdram_we_n                      (DRAM_WE_N),                     //                     .we_n
			// .sdram_clk_clk                   (DRAM_CLK),                   	//            sdram_clk.clk

			// HPS DDR3 SDRAM interface 
			// .hps_sdram_address				 (hps_sdram_address),
			// .hps_sdram_burstcount			 (8'b1),	
			// .hps_sdram_waitrequest			 (hps_sdram_waitrequest),	
			// .hps_sdram_writedata			 (hps_sdram_writedata),	
			// .hps_sdram_byteenable			 ({4{1'b1}}),	
			// .hps_sdram_write				 (hps_sdram_write),                   
			// .hps_sdram_readdata 			 (hps_sdram_readdata),                //                        .readdata
			// .hps_sdram_readdatavalid 		 (hps_sdram_readdatavalid),           //                        .readdatavalid
			// .hps_sdram_read 				 (hps_sdram_read),                    //  

			// Parallel Port
			.vid_pp_out_export 				 	(cmd_from_hps),

			// Clock Bridge
			.clock_bridge_0_in_clk_clk			(GPIO_1[1]),

			// FPGA to HPS FIFO
			.fifo_fpga_to_hps_in_writedata      (fpga_to_hps_in_writedata),      // fifo_fpga_to_hps_in.writedata
			.fifo_fpga_to_hps_in_write          (fpga_to_hps_in_write),          //                     .write
			.fifo_fpga_to_hps_in_csr_address    (32'd1), //(fpga_to_hps_in_csr_address),    //  fifo_fpga_to_hps_in_csr.address
			.fifo_fpga_to_hps_in_csr_read       (1'b1), //(fpga_to_hps_in_csr_read),       //                         .read
			.fifo_fpga_to_hps_in_csr_writedata  (),  //                         .writedata
			.fifo_fpga_to_hps_in_csr_write      (1'b0),      //                         .write
			.fifo_fpga_to_hps_in_csr_readdata   (fpga_to_hps_in_csr_readdata),    //                         .readdata
	
			// onchip SRAM
			// .onchip_sram_s1_address               (sram_address),               
			// .onchip_sram_s1_clken                 (sram_clken),                 
			// .onchip_sram_s1_chipselect            (sram_chipselect),            
			// .onchip_sram_s1_write                 (1'b0),                 
			// .onchip_sram_s1_readdata              (sram_readdata),              
			// .onchip_sram_s1_writedata             (sram_writedata),             
			// .onchip_sram_s1_byteenable            (4'b1111), 

			// mipi clock pll
			// .mipi_clock_sdram_clk_clk 			  (GPIO_1[1]),
			// .mipi_clock_ref_reset_reset 		  (0),

			// off chip sdram
			.sdram_s1_address				 	  (oc_sdram_address),
			.sdram_s1_byteenable_n			 	  ({4{1'b0}}),	
			.sdram_s1_chipselect 				  (1'b1),
			.sdram_s1_writedata			 	 	  (oc_sdram_writedata),	         //                        .readdatavalid
			.sdram_s1_read_n 				 	  (~oc_sdram_read),  
			.sdram_s1_write_n				 	  (~oc_sdram_write),                   
			.sdram_s1_readdata 			 	 	  (oc_sdram_readdata),                //                        .readdata
			.sdram_s1_readdatavalid 		 	  (oc_sdram_readdatavalid), 
			.sdram_s1_waitrequest			 	  (oc_sdram_waitrequest),	 

			// mipi clock pll
			// .mipi_clock_ref_clk_clk 		 	  (GPIO_1[1]),
			
//			.slider_switches_export          (SW),          						//      slider_switches.export
			.system_pll_ref_clk_clk          (CLOCK_50),          				//   system_pll_ref_clk.clk
			.system_pll_ref_reset_reset      (0)       								// system_pll_ref_reset.reset

		);


		///////////////////////////////////////////////////////////////////////////////////////////////
		// Instantiate an instance of the graphics and video controller circuit drawn as a schematic
		///////////////////////////////////////////////////////////////////////////////////////////////
			
		Graphics_and_Video_Controller		GraphicsController1 ( 
				.Reset_L							(RESET_L_WIRE),
				.Clock_50Mhz 					(CLOCK_50),
				.Address 						(IO_Address_WIRE),
				.DataIn 							(IO_Write_Data_WIRE),
				.DataOut 						(IO_Read_Data_WIRE),
				.IOEnable_L 					(IO_Enable_L_WIRE),
				.UpperByteSelect_L 			(IO_UpperByte_Select_L_WIRE),
				.LowerByteSelect_L 			(IO_LowerByte_Select_L_WIRE),
				.WriteEnable_L 				(IO_RW_WIRE),
				.GraphicsCS_L 					(IO_Enable_L_WIRE),
				
				.VGA_CLK						(VGA_CLK),
				.VGA_B 						(VGA_B),
				.VGA_G 						(VGA_G),
				.VGA_R							(VGA_R),
				.VGA_HS 						(VGA_HS),
				.VGA_VS						(VGA_VS),
				.VGA_BLANK_N 					(VGA_BLANK_N)

		 );
		
	
		///////////////////////////////////////////////////////////////////////////////////////////////
		// create an instance of the IO port with serial ports
		///////////////////////////////////////////////////////////////////////////////////////////////

		 OnChipSerialIO     SerialIOPorts (
				 
				 // Bridge Signals connecting to this component
				 
				 .Reset_L 						(RESET_L_WIRE),
				 .Clock_50Mhz 					(CLOCK_50),
				 .Address 						(IO_Address_WIRE),
				 .DataIn 						(IO_Write_Data_WIRE[7:0]),
				 .DataOut 						(IO_Read_Data_WIRE[7:0]),
				 .IOSelect_H 					(IO_Bus_Enable_WIRE),
				 .ByteSelect_L 				(IO_LowerByte_Select_L_WIRE),
				 .WE_L 							(IO_RW_WIRE),
				 .IRQ_H 							(IO_IRQ_WIRE),
				 
				 // Real World Signals brought out to Header connections
				 
				 .RS232_RxData					(GPIO_0[29]),
				 .RS232_TxData					(GPIO_0[27]),

				 .GPS_RxData 					(GPIO_0[28]),
				 .GPS_TxData 					(GPIO_0[26]),

				 .BlueTooth_RxData 			(GPIO_0[32]),
				 .BlueTooth_TxData 			(GPIO_0[34]),
				 
				 .TouchScreen_RxData 		(GPIO_0[11]),
				 .TouchScreen_TxData 		(GPIO_0[10])
		);

		//=======================================================
		// Controls for Qsys sram slave exported in system module
		//=======================================================
		wire [31:0] sram_readdata ;
		reg [31:0] sram_writedata ;
		reg [7:0] sram_address; 
		wire sram_clken = 1'b1;
		wire sram_chipselect = 1'b1;
		reg [7:0] state ;

		//=======================================================
		// Controls for Qsys SDRAM controller exported in system module
		//=======================================================
		// wire [24:0] 	off_chip_sdram_address;
		// wire [1:0] 		off_chip_sdram_byteenable_n;
		// wire  			off_chip_sdram_chipselect;
		// wire [31:0] 	off_chip_sdram_writedata;
		// wire  			off_chip_sdram_read_n;
		// wire 			off_chip_sdram_write_n;
		// wire [31:0] 	off_chip_sdram_readdata;
		// wire  			off_chip_sdram_readdatavalid;
		// wire  			off_chip_sdram_waitrequest;

		//=======================================================
		// Controls for FPGA_to_HPS FIFO
		//=======================================================

		reg[31:0] fpga_to_hps_in_csr_readdata ;
		reg fpga_to_hps_in_csr_read ; // status regs read cmd
		reg [7:0] FPGA_to_HPS_state ;

		wire [31:0] fpga_to_hps_in_writedata ; 
		wire fpga_to_hps_in_write ; // write command
		wire [31:0] fpga_to_hps_in_csr_address = 32'd1 ; // fill_level

		assign fpga_to_hps_in_write = FPGA_to_HPS_state == 5 ? 1'b1 : 1'b0;
		assign fpga_to_hps_in_writedata = {RED, GREEN, BLUE}; 

		//=======================================================
		// Controls for HPS SDRAM interface
		//=======================================================

		// assign hps_sdram_write = FPGA_to_HPS_state == 1 ? 1'b1 : 1'b0;
		// assign hps_sdram_read = FPGA_to_HPS_state == 2 ? 1'b1 : 1'b0;
		// assign hps_sdram_address = (FPGA_to_HPS_state == 2 ? SDRAM_counter2 : SDRAM_counter1);
		// assign hps_sdram_writedata = {6'b0, rgb_out};

		wire [24:0] oc_sdram_address;
		wire [15:0] oc_sdram_writedata, oc_sdram_readdata;
		wire oc_sdram_read, oc_sdram_write, oc_sdram_readdatavalid, oc_sdram_waitrequest;

		wire [11:0] pixel_out;
		wire pixel_valid;

		reg [15:0] sdram_out;

		always @(posedge CLOCK_50) begin
			if (~fpga_to_hps_fifo_rst_n) begin
				sdram_out <= 0;
			end else if (oc_sdram_readdatavalid) begin
				sdram_out <= oc_sdram_readdata;
			end
		end

		assign oc_sdram_write = FPGA_to_HPS_state == 1 ? pixel_valid & ~oc_sdram_waitrequest : 1'b0;
		assign oc_sdram_read = FPGA_to_HPS_state == 2 ? ~f2h_fifo_full : 1'b0;
		assign oc_sdram_address = (FPGA_to_HPS_state == 1 ? SDRAM_counter1 : SDRAM_counter2);
		assign oc_sdram_writedata = {4'b0, pixel_out};

		wire MIPI_PIXEL_VS, MIPI_PIXEL_HS;
		assign MIPI_PIXEL_VS = GPIO_1[20];
		assign MIPI_PIXEL_HS = GPIO_1[22];

		wire [9:0] OUT_MIPI_PIXEL_D;
		wire OUT_MIPI_PIXEL_VS, OUT_MIPI_PIXEL_HS;
		wire [8:0] RED, GREEN, BLUE;

		assign OUT_MIPI_PIXEL_D =  sdram_out[9:0];
		assign OUT_MIPI_PIXEL_HS = sdram_out[10];
		assign OUT_MIPI_PIXEL_VS = sdram_out[11];
		// assign OUT_MIPI_PIXEL_HS = Width_counter == VIDEO_W;
		// assign OUT_MIPI_PIXEL_VS = Height_counter == VIDEO_H || (Width_counter == 0 && Height_counter == 0);

		
		//------ CMOS CCD_DATA TO RGB_DATA -- 
		RAW2RGB_J				u4	(	
			.RST          ( OUT_MIPI_PIXEL_VS ),
			.iDATA        ( OUT_MIPI_PIXEL_D ),		
			//-----------------------------------
			.VGA_CLK      ( CLOCK_50 ),
			.READ_Request ( 1'b1 ),
			.VGA_VS       ( OUT_MIPI_PIXEL_VS ),	
			.VGA_HS       ( OUT_MIPI_PIXEL_HS ), 

			.oRed         ( RED  ),
			.oGreen       ( GREEN),
			.oBlue        ( BLUE )
		);

		//=======================================================
		// Controls for Camera RGB to SDRAM
		//=======================================================
		wire f2h_fifo_full;
		assign f2h_fifo_full = fpga_to_hps_in_csr_readdata[0];
		
		wire fpga_to_hps_fifo_rst_n;
		assign fpga_to_hps_fifo_rst_n = KEY[0];

		wire output_finished;
		wire transfer_finished;

		// assign save_frame = FPGA_to_HPS_state == 1;

		assign output_finished = SDRAM_counter1 == 32'd307200;
		assign transfer_finished = SDRAM_counter2 == 32'd307200;
		assign start_transmission = cmd_from_hps[0]; 

		reg save_frame;
		always @(posedge GPIO_1[1]) begin
			if (~fpga_to_hps_fifo_rst_n) begin
				save_frame <= 0;
			end else if (output_finished) begin
				save_frame <= 0;
			end else if (MIPI_PIXEL_VS & MIPI_PIXEL_HS) begin
				save_frame <= cmd_from_hps[0];
			end
		end

		always @(posedge CLOCK_50) begin 
			// reset state machine and read/write controls
			if (~fpga_to_hps_fifo_rst_n) begin
				FPGA_to_HPS_state <= 8'd0 ;
			end

			//=======================================================
			// State 0: Waiting for Start
			//=======================================================
			if (FPGA_to_HPS_state==0) begin
				FPGA_to_HPS_state <= start_transmission ? 8'd1 : 8'd0;
			end

			//=======================================================
			// State 1: Saving Frame in SDRAM
			//=======================================================
			if (FPGA_to_HPS_state==1) begin
				FPGA_to_HPS_state <= output_finished ? 8'd2 : 8'd1;
			end

			//=======================================================
			// State 2: Sending Data From SDRAM to HPS
			//=======================================================
			if (FPGA_to_HPS_state==2) begin // read from sdram
				FPGA_to_HPS_state <= oc_sdram_read ? 8'd3 : 8'd2;
			end

			if (FPGA_to_HPS_state==3) begin // wait for readdatavalid
				FPGA_to_HPS_state <= oc_sdram_readdatavalid ? 8'd4 : 8'd3;
			end

			if (FPGA_to_HPS_state==4) begin // wait for RAW_2_RGB Model and HPS fifo not full
				FPGA_to_HPS_state <= f2h_fifo_full ? 8'd4 : 8'd5;
			end

			if (FPGA_to_HPS_state==5) begin // send to hps
				FPGA_to_HPS_state <= transfer_finished ? 8'd0 : 8'd2;
			end
		end

		assign LEDR = {FPGA_to_HPS_state[2:0], 4'h0, transfer_finished, output_finished, start_transmission};

		//=======================================================
		// Addresses
		//=======================================================
		reg [32:0] SDRAM_counter1, SDRAM_counter2;

		always @(posedge CLOCK_50) begin
			if (~fpga_to_hps_fifo_rst_n) begin
				SDRAM_counter1 <= 0;
			end else if (FPGA_to_HPS_state==1) begin
				SDRAM_counter1 <= SDRAM_counter1 + oc_sdram_write;
			end else begin
				SDRAM_counter1 <= 0;
			end
		end

		always @(posedge CLOCK_50) begin
			if (~fpga_to_hps_fifo_rst_n) begin
				SDRAM_counter2 <= 0;
			end else if (FPGA_to_HPS_state==4) begin
				SDRAM_counter2 <= SDRAM_counter2 + ~f2h_fifo_full;
			end else if (FPGA_to_HPS_state==0) begin
				SDRAM_counter2 <= 0;
			end
		end

		parameter VIDEO_W	= 640;
		parameter VIDEO_H	= 480;

		reg [32:0] Width_counter, Height_counter;

		always @(posedge CLOCK_50) begin
			if (~fpga_to_hps_fifo_rst_n) begin
				Width_counter <= 0;
				Height_counter <= 0;
			end else if (FPGA_to_HPS_state==4) begin
				if (Width_counter == VIDEO_W && fpga_to_hps_in_write) begin
					Width_counter <= 0;
					Height_counter <= Height_counter + 1;
				end else begin
					Width_counter <= Width_counter + fpga_to_hps_in_write;
					Height_counter <= Height_counter;
				end
			end else begin
				Width_counter <= 0;
				Height_counter <= 0;
			end
		end


		///////////////////////////////////////////////////////////////////////////////////////////////
		// create an instance of the D8M camera
		///////////////////////////////////////////////////////////////////////////////////////////////
		
		Camera D8M_Camera (
			//////////// CLOCK //////////
			.CLOCK_50 					(CLOCK_50),
			.CLOCK2_50 					(CLOCK2_50),
			.CLOCK3_50 					(CLOCK3_50),

			//////////// MIPI CAMERA (D8M) //////////
			.CAMERA_I2C_SCL				(GPIO_1[26]),	
			.CAMERA_I2C_SDA				(GPIO_1[27]),	
			.CAMERA_PWDN_n				(GPIO_1[25]),	
			.MIPI_CS_n					(GPIO_1[23]),
			.MIPI_I2C_SCL				(GPIO_1[30]),	
			.MIPI_I2C_SDA				(GPIO_1[31]),	
			.MIPI_MCLK					(GPIO_1[28]),
			.MIPI_PIXEL_CLK				(GPIO_1[1]),	
			.MIPI_PIXEL_D				(GPIO_1[12:3]),	
			.MIPI_PIXEL_HS				(GPIO_1[22]),	
			.MIPI_PIXEL_VS				(GPIO_1[20]),	
			.MIPI_REFCLK				(GPIO_1[18]),	
			.MIPI_RESET_n				(GPIO_1[24]),	
			
			.KEY 						(KEY),
			.SW 						(SW),
			.pixel_out 					(pixel_out),
			.pixel_valid  				(pixel_valid),
			.waitreq 					(oc_sdram_waitrequest),
			.save_frame 				(save_frame)

			// SDRAM interface
			
			// .DRAM_ADDR                      (DRAM_ADDR),                     //                sdram.addr
			// .DRAM_BA                       	(DRAM_BA),                       //                     .ba
			// .DRAM_CAS_N                     (DRAM_CAS_N),                    //                     .cas_n
			// .DRAM_CKE                       (DRAM_CKE),                      //                     .cke
			// .DRAM_CS_N                      (DRAM_CS_N),                     //                     .cs_n
			// .DRAM_DQ                       	(DRAM_DQ),                       //                     .dq
			// .Temp_SDRAM_DQM 				(Temp_SDRAM_DQM),                //                     .dqm
			// .DRAM_RAS_N                     (DRAM_RAS_N),                    //                     .ras_n
			// .DRAM_WE_N                      (DRAM_WE_N),                     //                     .we_n
			// .DRAM_CLK                   	(DRAM_CLK)                   	// 
			
		);

		HEX_DISPLAY addr_display (
			// .wraddr		({fpga_to_hps_in_write, 3'h0, f2h_fifo_full, 3'h0, cmd_from_hps[0], 3'h0, output_finished, 3'h0, FPGA_to_HPS_state[0]}),
			.wraddr 	(oc_sdram_address),
			.HEX0 		(HEX0),
			.HEX1 		(HEX1),
			.HEX2 		(HEX2),
			.HEX3 		(HEX3),
			.HEX4 		(HEX4),
			.HEX5 		(HEX5)
		);

		// Map 16 bit memory upper and lower data byte strobes to individual wires
		assign RESET_L_WIRE 	= 1'b1;	 
		
		// connections to wires on the top level to invert signals coming from the bridge
		
		assign IO_Enable_L_WIRE 				= ~IO_Bus_Enable_WIRE;
		assign IO_UpperByte_Select_L_WIRE 	= ~IO_Byte_Enable_WIRE[1];		
		assign IO_LowerByte_Select_L_WIRE 	= ~IO_Byte_Enable_WIRE[0];	
	
		// process to generate an acknowledge for the IO Bridge 1 clock cycle after bridge IO BUS ENABLE and then remove it 
		always@(posedge CLOCK_50)
		begin
			IO_ACK_WIRE <= IO_Bus_Enable_WIRE;
		end
endmodule